---------------------------------------------------------------------------------------------------
--
-- Title       : Frequency Divider
-- Design      : WORK
-- Author      : ManRares
-- Company     : UT Cluj-Napoca
--
---------------------------------------------------------------------------------------------------
--
-- File        : Frequency
-- Generated   : Fri Apr 17 18:27:28 2020
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------