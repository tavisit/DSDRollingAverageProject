---------------------------------------------------------------------------------------------------
--
-- Title       : Data_Generator
-- Design      : WORK
-- Author      : Man Rares
-- Company     : UT Cluj-Napoca
--
---------------------------------------------------------------------------------------------------
--
-- File        : Data_Generator.vhd
-- Generated   : Tue Apr 28 13:57:05 2020
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity Data_Generator is
	port ( Reset: in std_logic;
		   Control: in std_logic_vector(2 downto 0);
		   SystemClock: in std_logic;
		   Data: out std_logic_vector(7 downto 0);
		   DataClock: inout std_logic);
end Data_Generator;

architecture DataGen of Data_Generator is
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- 													                       Necessary components																							  --
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	component FrequencyDivider is
		port (SysClk, Reset: in std_logic;
	      DataClk: out std_logic);	   
	end component;
	
	component SquareWave is
		port (ClkIn, Reset, enable: in std_logic;
		  	  ClkOut: inout std_logic;
		  	  DataOut: out std_logic_vector (7 downto 0));	   
	end component;
	
	component Mux_8 is	
	PORT ( A: in Std_logic_vector(7 downto 0);
		   B : in Std_logic_vector(7 downto 0);
		   C : in Std_logic_vector(7 downto 0);
		   D : in Std_logic_vector(7 downto 0);
		   E : in Std_logic_vector(7 downto 0);
		   F : in Std_logic_vector(7 downto 0);
		   G : in Std_logic_vector(7 downto 0);
		   H : in Std_logic_vector(7 downto 0);
		   Sel: in Std_logic_vector(2 downto 0);
		   Data : out Std_logic_vector(7 downto 0));
	end component;
															  	
	component Pseudo0_15 is
  		port ( cout:out std_logic_vector (7 downto 0);
   		 	   enable, clk, reset :in  std_logic);
	end component;
	
	component Pseudo0_255 is
  		port ( cout:out std_logic_vector (7 downto 0);
   		 	   enable, clk, reset :in  std_logic);                
	end component;
	
	component Reg is
		port ( Clk: in std_logic;
		   	   D: in std_logic_vector(7 downto 0);
		   	   Q: out std_logic_vector(7 downto 0));
	end component;
	
	component SixDigit1 is
  		port ( cout:out std_logic_vector (7 downto 0);
   		       enable, clk, reset :in  std_logic);
	end component;
	
	component SixDigit2 is
  		port ( cout:out std_logic_vector (7 downto 0);
   		 	   enable, clk, reset :in  std_logic);
	end component;
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- 													                      End of Necessary components																					  --		  
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- 													                       Necessary SIGNALS																							  --
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
							   
	signal SqWvClk: std_logic;
	signal DaClk: std_logic;
	signal A: std_logic_vector(7 downto 0);
	signal B: std_logic_vector(7 downto 0);
	signal C: std_logic_vector(7 downto 0);
	signal D: std_logic_vector(7 downto 0);
	signal E: std_logic_vector(7 downto 0);
	signal DataAux: std_logic_vector(7 downto 0);
	
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- 													                      End of Necessary SIGNALS																						  --
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
begin

		FreqDiv: FrequencyDivider Port Map(SystemClock, Reset, DaClk);

			SqWv: SquareWave Port Map(DaClk, Reset, '1', SqWvClk, A);
			SD1: SixDigit1 Port Map(B, '1', DaClk, Reset);
			SD2: SixDigit2 Port Map(C, '1', DaClk, Reset);
			PRNG1: Pseudo0_15 Port Map(D, '1', DaClk, Reset);
			PRNG2: Pseudo0_255 Port Map(E, '1', DaClk, Reset);
			MUXData: MUX_8 Port Map("00000000", A, B, C, "00000000", "00000000", E, "00000000", Control, DataAux);
			MUXClock: MUX_8 Port Map(DaClk, SqWvClk, DaClk, DaClk, DaClk, DaClk, DaClk, DaClk, Control, DataClock);
			Regi: Reg Port Map(DataClock, DataAux, Data);
		
end DataGen;		