---------------------------------------------------------------------------------------------------
--
-- Title       : Filter
-- Design      : Project
-- Author      : OctavianMatei
-- Company     : UT Cluj-Napoca
--
---------------------------------------------------------------------------------------------------
--
-- File        : Filter.vhd
-- Generated   : Sun Apr 12 16:46:40 2020
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {Filter} architecture {Filter}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Filter is
	PORT(RESET,DATA_CLOCK : IN STD_LOGIC;
		DATA : IN STD_LOGIC_VECTOR(7 downto 0);	  
		Length: IN STD_LOGIC_VECTOR(2 downto 0);
		OUTPUT: OUT STD_LOGIC_VECTOR(7 downto 0));
end Filter;

--}} End of automatically maintained section

architecture Filter of Filter is  
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- 													                       Necessary components																							  --
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
component MainRegister is 
	PORT(RESET,CLK : IN STD_LOGIC;
	DATA : IN STD_LOGIC_VECTOR(7 downto 0);       --The Input data
	OUTPUT : INOUT STD_LOGIC_VECTOR(127 downto 0)); -- The Output stores every one of the 8 bit numbers, 16 in total
end component;

component MUX is	
	PORT ( A: IN STD_LOGIC_VECTOR(8 downto 0);
	B : IN STD_LOGIC_VECTOR(9 downto 0);
	C : IN STD_LOGIC_VECTOR(10 downto 0);
	D : IN STD_LOGIC_VECTOR(11 downto 0);
	SELECTION_LENGTH: IN STD_LOGIC_VECTOR(2 downto 0);
	SUM : OUT STD_LOGIC_VECTOR(11 downto 0));
end component;

component HexConverter is
	PORT( 	CLK : IN STD_LOGIC;
			INPUT:IN STD_LOGIC_VECTOR(7 downto 0 );	--INPUT SEGMENTED IN TWO PARTS
		  OUTPUT1,OUTPUT2: OUT STD_LOGIC_VECTOR(6 downto 0));
end component;
--lENGTH CONTROLS HOW MUCH TO SHIFT
--SHIFT LENGTH(1 DOWNTO 0)
component ShiftRegister is
	port(
	D: in STD_LOGIC_vector(11 downto 0);
	Length : IN STD_LOGIC_VECTOR (2 downto 0);
	     clock, RESET: in STD_LOGIC;
		 q: inout STD_LOGIC_vector(11 downto 0));
end component;
--NBITADDER
--WILL BE USED WITH NUMBEROFINPUTS AS FOLLOWS:
--8 FOR THE FIRST LAYER
--9 FOR THE SECOND
--10 FOR THE THIRD
--11 FOR THE FOURTH
component NBitAdder is	
  generic(
        numberOfInputs : Integer := 8
    ); port(
        cin     : in std_logic;
        inputs1 : in std_logic_vector(numberOfInputs-1 downto 0);
        inputs2 : in std_logic_vector(numberOfInputs-1 downto 0);
        outputs : out std_logic_vector(numberOfInputs downto 0)
    );
end component;	 
SIGNAL OUTPUTSMALL : STD_LOGIC_VECTOR(5 downto 0);
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- 													                       Necessary components																							  --
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
begin

end Filter;
